module or ();