module and (
    
);
