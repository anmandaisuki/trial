module or (
    input logic a ;
    output logic b;
    input logic c;

);