module or (
    input logic a ;
    output logic b;

);